----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 21.11.2015 16:58:00
-- Design Name: 
-- Module Name: comp - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity comp is
    Port ( CLOCK    : in STD_LOGIC                    ;
           RPS      : in STD_LOGIC_VECTOR (7 downto 0);
           SETPOINT : in STD_LOGIC_VECTOR (7 downto 0);
           RES      : out STD_LOGIC_VECTOR(7 downto 0);
           POS      : out STD_LOGIC                  );
end comp;

architecture Behavioral of comp is
    signal result : std_logic_vector(7 downto 0);
    signal rot    : std_logic_vector(7 downto 0);
    signal sp     : std_logic_vector(7 downto 0);
begin

RES<=result   ;
rot<=RPS      ;
sp <=SETPOINT ;

process(rot,sp,CLOCK)
begin
    if rising_edge(CLOCK) then
        if(SETPOINT>=RPS) then
            result<=std_logic_vector(unsigned(sp)-unsigned(rot));
            POS   <='1';
        else
            result<=std_logic_vector(unsigned(rot)-unsigned(sp));
            POS   <='0';
        end if;
    end if;
end process;


end Behavioral;
